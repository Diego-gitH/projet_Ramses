library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ramses is port(
	clock0 : in std_logic;
	clock1 : in std_logic;
	buttons : in std_logic_vector(0 to 3) := "000";
	first_7segment : out std_logic_vector(3 downto 0);
	second_7segment : out std_logic_vector(3 downto 0);
	rows_matrix : out std_logic_vector(0 to 6);
	cols_matrix : out std_logic_vector(0 to 4);
	reset : in std.logic;
);
end entity ramses;

architecture Behavioral of ramses is
	constant ROWS : integer := 7;
	constant COLS : integer := 5;
	
begin
	
	
end architecture Behavioral;